wire [99:0] my_vector;
assign out = my_vector[10]