module start (
    output zero;
);

    assign zero = 0;
    
endmodule