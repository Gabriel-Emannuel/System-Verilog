// module top_module ( input a, input b, output out );
//     mod_a manager(.out(out), .in1(a), .in2(b));
// endmodule

// module top_module ( input a, input b, output out );
//     mod_a manager(a, b,out);
// endmodule